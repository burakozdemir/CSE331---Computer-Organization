module ALU_testbench();

reg [3:0] ALUcontrol;
reg [31:0] A,B;
wire [31:0] ALUout;
wire zero;

ALU x(ALUcontrol,A,B,ALUout,zero);

initial begin
ALUcontrol = 4'b1000 ;//a + b
A = 32'b00000000010000100101000000100000; 
B = 32'b00000000010000100101000000100000; #10;
ALUcontrol = 4'b1100 ;//a & b
A = 32'b00000000010000100101000000100000; 
B = 32'b00000000010000100101000000100000; #10;
ALUcontrol = 4'b1001 ;//a - b
A = 32'b00000000010000100101000000100000; 
B = 32'b00000000010000100101000000100000; #10;
ALUcontrol = 4'b0100 ;//a or b
A = 32'b11111111111111111111111111100000; 
B = 32'b00000000010000100101000000100000; #10;
ALUcontrol = 4'b1011 ;//b << 1
A = 32'b00000000000000000000000000000111; 
B = 32'b00000000000000000000000000001110; #10;
ALUcontrol = 4'b1010 ;//b >> 1
A = 32'b00000000000000000000000000000111; 
B = 32'b00000000000000000000000000001110; #10;
ALUcontrol = 4'b0010 ;//b >>> 1
A = 32'b00000000000000000000000000000111; 
B = 32'b00000000000000000000000000001110; #10;
ALUcontrol = 4'b111 ;//rd = 1 or 0
A = 32'b00000000000000000000000000000111; 
B = 32'b00000000000000000000000000001110; #10;

end

initial begin
  $monitor("Test-Time:%2d, ALUcntrl: %4b ,A: %32b,B: %32b,Result: %32b",
            $time,ALUcontrol,A,B,ALUout);
end

endmodule